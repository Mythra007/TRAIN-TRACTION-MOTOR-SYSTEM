* Final Complete Train Traction System Simulation - Version 29 (Arithmetic Logic Final)

.title Lam Research Train Traction System System - Final Submission V29
.save all
.probe alli

* --- Model Definitions ---
.model D_GENERIC D(Is=1n Rs=0.1) ; Generic Diode model

* --- Model Definitions ---
.model __D1 D(Is=1n Rs=0.1) ; Diode model from KiCAD netlist
.model __D2 D(Is=1n Rs=0.1) ; Diode model from KiCAD netlist


.model __Q1 VDMOS(Vto=1 Kp=50m Rd=0.01 Rs=0.01) ; Model for KiCAD Q1 (Main Buck Switch)
.model __Q2 VDMOS(Vto=1 Kp=50m Rd=0.01 Rs=0.01) ; Model for KiCAD Q2 (Motor Branch Switch)
.model __Q3 VDMOS(Vto=1 Kp=50m Rd=0.01 Rs=0.01) ; Model for KiCAD Q3 (Regeneration Switch)
.model M_BRAKE_VDMOS VDMOS(Vto=1 Kp=50m Rd=0.01 Rs=0.01) ; Model for Braking Resistor Switch

* --- Global Parameters (for easier tuning) ---
.param PWM_FREQ = 100k
.param PWM_PERIOD = {1/PWM_FREQ}
.param PWM_ON_MAX = 5 ; Max voltage for PWM ON state (e.g., 5V for IGBT gate)
.param PID_MAX_OUT = 5 ; Max output voltage of PID controller (maps to PWM_ON_MAX)

.param R_SENSE_VAL = 0.01 ; KiCAD R2 value (Motor current sense shunt)
.param R_MOTOR_RA_VAL = 0.5 ; KiCAD R3 value (Motor Armature Resistance)
.param L_MOTOR_LA_VAL = 10m ; KiCAD L2 value (Motor Armature Inductance)
.param K_EMF = 0.05 ; Back EMF constant (V/(rad/s))

.param CURRENT_THRESHOLD_V = 0.15 ; Op-amp threshold for overcurrent (V)
.param STALL_CURRENT_THRESHOLD_V = 0.05 ; Op-amp threshold for stall current (V)
.param STALL_SPEED_THRESHOLD_V = 0.5 ; Op-amp threshold for stall speed (V)
.param TEMP_THRESHOLD_V = 80 ; Op-amp threshold for overtemperature (V)
.param INSULATION_FAULT_THRESHOLD_V = 0.2 ; Threshold for insulation health (normalized 0-1)
.param STUCK_DURATION_THRESHOLD_S = 10u ; Time for PWM/Sensor stuck fault detection (s)

.param REGEN_CAP_VAL = 100m ; Value for main regenerative capacitor (Farads)
.param BRAKE_RESISTOR_VAL = 5 ; Value for braking resistor (Ohms)
.param L_REGEN_VAL = 1m ; Regenerative Inductor (Henrys)

.param TEG_GAIN_VAL = 0.05

.param VCC_LIMIT = 5 ; Matches VCC_RAIL voltage
.param VEE_LIMIT = -5 ; Matches VEE_RAIL voltage

.param C_IN_VAL = 100u ; Value for KiCAD C4 (Input Capacitor)
.param C_BUCK_OUT_VAL = 470u ; Value for Buck Output Capacitor (explicitly added)
.param L_BUCK_VAL = 100u ; Value for KiCAD L1 (Buck Inductor)

.param RPULLDOWN = 1Meg ; Value for pull-down resistors on behavioral outputs

* --- Power Supplies ---
VCC_RAIL VCC GND DC 5V
VEE_RAIL VEE GND DC -5V

* --- Ideal Op-Amp Subcircuit ---
.subckt IDEAL_OPAMP_SUB NON_INV_IN INV_IN OUT_NODE
E_gain_output Output_unclamped GND VALUE={(V(NON_INV_IN) - V(INV_IN)) * 1e5}
E_clamped_output OUT_NODE Output_unclamped VALUE={LIMIT(V(Output_unclamped), VEE_LIMIT, VCC_LIMIT)}
.ends IDEAL_OPAMP_SUB

* --- PID Controller Subcircuit ---
.subckt PID_CONTROLLER VREF VACTUAL_SPEED VPID_OUT GND_NODE
.param Kp_val = 10
.param Ki_val = 100
.param Kd_val = 0.01
E_error ERROR_NODE GND_NODE VALUE = {V(VREF) - V(VACTUAL_SPEED)}
E_P P_TERM GND_NODE VALUE = {Kp_val * V(ERROR_NODE)}
C_int INTEGRAL_NODE GND_NODE 1uF
R_int_feedback ERROR_NODE INTEGRAL_NODE 1meg
E_I I_TERM GND_NODE VALUE = {Ki_val * V(INTEGRAL_NODE)}
R_deriv_input ERROR_NODE DERIV_NODE 1k
C_deriv_shunt DERIV_NODE GND_NODE 1nF
E_D D_TERM GND_NODE VALUE = {Kd_val * ddt(V(ERROR_NODE))}
E_PID_OUT VPID_OUT GND_NODE VALUE = {V(P_TERM) + V(I_TERM) + V(D_TERM)}
.ends PID_CONTROLLER

* --- Main Circuit Netlist ---

* --- Threshold Voltage Sources ---
V4_src /CURRENT_THRESHHOLD GND DC {CURRENT_THRESHOLD_V}
V9_src /STALL_CURRENT_THRESHHOLD GND DC {STALL_CURRENT_THRESHOLD_V}
V10_src /STALL_SPEED_THRESHHOLD GND DC {STALL_SPEED_THRESHOLD_V}
V5_src /TEMP_THRESHHOLD GND DC {TEMP_THRESHOLD_V}
V_INSULATION_THRESHOLD INSULATION_THRESHOLD_NODE GND DC {INSULATION_FAULT_THRESHOLD_V}
V29_src /USER_CONTROLLED_BRAKE GND DC 0V
R_USER_CTRL_BRAKE_PULLDOWN /USER_CONTROLLED_BRAKE GND {RPULLDOWN}

* --- Reference Inputs ---
V3 /V_REF GND PWL(0 0 1s 50 5s 80 8s 50 10s 0)

* --- Input Stage (KiCAD V1, C4) ---
V1_source V_INPUT_MAIN GND DC 100V ; KiCAD V1: Main DC Input Voltage Source
C4_INPUT V_INPUT_MAIN GND {C_IN_VAL} ; KiCAD C4: Input Filter Capacitor, across source and GND

* --- Buck Converter (KiCAD Q1, L1, D1, C_BUCK_OUTPUT_FILTER) ---
* Q1 from your schematic is the main buck switch.
M1_BUCK_MAIN V_INPUT_MAIN PWM_OUT_NODE L1_INPUT_NODE L1_INPUT_NODE __Q1 ; KiCAD Q1: Main Buck Switch (Drain=V_INPUT_MAIN, Gate=PWM_OUT_NODE, Source=L1_INPUT_NODE)
L1_BUCK L1_INPUT_NODE BUCK_OUTPUT_NODE {L_BUCK_VAL} ; KiCAD L1: Buck Inductor
D1_FREEWHEELING GND BUCK_OUTPUT_NODE D_GENERIC ; KiCAD D1: Freewheeling Diode (Anode=GND, Cathode=BUCK_OUTPUT_NODE)
C_BUCK_OUTPUT_FILTER BUCK_OUTPUT_NODE GND {C_BUCK_OUT_VAL} ; Buck Output Filter Capacitor
R_CBUCK_SHUNT BUCK_OUTPUT_NODE GND 1G ; Shunt across output capacitor for DC stability

* --- Motor Branch (KiCAD Q2, R2, R3, L2, E1) ---
* Q2 from your schematic is the motor branch switch.
M2_MOTOR_BRANCH_SWITCH BUCK_OUTPUT_NODE Q2_GATE_NODE MOTOR_ARMATURE_INPUT MOTOR_ARMATURE_INPUT __Q2 ; KiCAD Q2: Motor Branch Switch
* Control for Q2 (always ON for normal operation, or controlled if needed)
V_Q2_CTRL Q2_GATE_NODE GND DC 5V ; Always ON (5V for gate)
R_Q2_GATE_SERIES Q2_GATE_SOURCE_NODE Q2_GATE_NODE 100u

R2_MOTOR_SENSE_SHUNT MOTOR_ARMATURE_INPUT MOTOR_RA_LA_NODE {R_SENSE_VAL} ; KiCAD R2: Motor current sense shunt
R3_MOTOR_ARMATURE_RES MOTOR_RA_LA_NODE MOTOR_L_NODE {R_MOTOR_RA_VAL} ; KiCAD R3: Armature Resistance
L2_MOTOR_ARMATURE_IND MOTOR_L_NODE /MOTOR_SPEED_NODE {L_MOTOR_LA_VAL} ; KiCAD L2: Armature Inductance
E1_BACK_EMF /MOTOR_SPEED_NODE GND VALUE={K_EMF * V(/MOTOR_SPEED_NODE)} ; KiCAD E1: Back EMF
R_L_MOTOR_SHUNT L2_MOTOR_ARMATURE_IND MOTOR_L_NODE 1u ; Small series R for inductor DC stability

* --- Current Sense Amplifier (Behavioral - Replaced KiCAD U1) ---
* Now sensing across R2_MOTOR_SENSE_SHUNT. Note: V(MOTOR_ARMATURE_INPUT) is node before R2 (shunt), V(MOTOR_RA_LA_NODE) is node after R2.
E_CS_AMP_FINAL CURRENT_SENSE_OUT GND VALUE={MIN(MAX(0, (V(MOTOR_ARMATURE_INPUT) - V(MOTOR_RA_LA_NODE)) * 100), VCC_LIMIT)} ; Gain 100, clamped


* --- Motor Load (Behavioral - Arithmetic Logic) ---
G_load /MOTOR_SPEED_NODE GND VALUE = { (10 * V(/MOTOR_SPEED_NODE)) + (MAX(0.0, (time - 3s)) * MAX(0.0, (5s - time)) * 10 * V(/MOTOR_SPEED_NODE) / (2s*1s)) + (MAX(0.0, (time - 7s)) * MAX(0.0, (9s - time)) * 20 * V(/MOTOR_SPEED_NODE) / (2s*1s)) }


* --- PID Controller (Behavioral) ---
X_PID_CONTROLLER /V_REF /MOTOR_SPEED_NODE PID_OUT_NODE GND PID_CONTROLLER
R_PID_OUT_PULLDOWN PID_OUT_NODE GND {RPULLDOWN}

* --- PWM Generator (Behavioral - Arithmetic Logic) ---
E_PWM_GEN PWM_OUT_NODE GND VALUE = {(MAX(0.0, ( (V(PID_OUT_NODE) / PID_MAX_OUT * PWM_PERIOD) - (time - floor(time/PWM_PERIOD)*PWM_PERIOD) )) * PWM_ON_MAX) / (PWM_PERIOD)}


* --- Fault Detection System (Behavioral) ---
* All comparators replaced with basic E-sources that output 0 or 1.


* Overcurrent Fault (KiCAD U7 equivalent)
E_FAULT_OVERCURRENT FAULT_OVERCURRENT_FLAG GND VALUE={MIN(MAX(0.0, (V(CURRENT_SENSE_OUT) - V(/CURRENT_THRESHHOLD)))*1k, 1)}
R_OC_FLAG_PULLDOWN FAULT_OVERCURRENT_FLAG GND {RPULLDOWN}

* Motor Stall (KiCAD U8 & U9 equivalents)
E_FAULT_STALL_SPEED_LOW FAULT_STALL_SPEED_LOW_FLAG GND VALUE={MIN(MAX(0.0, (V(/STALL_SPEED_THRESHHOLD) - V(/MOTOR_SPEED_NODE)))*1k, 1)}
R_SS_FLAG_PULLDOWN FAULT_STALL_SPEED_LOW_FLAG GND {RPULLDOWN}
E_FAULT_STALL_CURRENT_HIGH STALL_CURRENT_HIGH_FLAG GND VALUE={MIN(MAX(0.0, (V(CURRENT_SENSE_OUT) - V(/STALL_CURRENT_THRESHHOLD)))*1k, 1)}
R_SC_FLAG_PULLDOWN STALL_CURRENT_HIGH_FLAG GND {RPULLDOWN}

E_COMBINED_FAULT_STALL FAULT_STALL_FLAG GND VALUE={V(FAULT_STALL_SPEED_LOW_FLAG) * V(STALL_CURRENT_HIGH_FLAG)} ; AND logic is multiplication
R_STALL_FLAG_PULLDOWN FAULT_STALL_FLAG GND {RPULLDOWN}

* PWM Stuck (Behavioral)
E_PWM_STUCK_COND_A PWM_STUCK_COND_A_NODE GND VALUE={MAX(0.0, (V(PID_OUT_NODE) - 4))} ; No *1k here, it's a condition flag
R_PWM_STUCK_COND_A_PULLDOWN PWM_STUCK_COND_A_NODE GND {RPULLDOWN}
E_PWM_STUCK_COND_B PWM_STUCK_COND_B_NODE GND VALUE={MAX(0.0, (1 - V(PWM_OUT_NODE)))} ; No *1k here, it's a condition flag
R_PWM_STUCK_COND_B_PULLDOWN PWM_STUCK_COND_B_NODE GND {RPULLDOWN}
E_PWM_STUCK_RAW PWM_STUCK_RAW_NODE GND VALUE={ MIN(1, V(PWM_STUCK_COND_A_NODE) * V(PWM_STUCK_COND_B_NODE)) } ; Combined AND, clamped to 1
R_PWM_STUCK_RAW_PULLDOWN PWM_STUCK_RAW_NODE GND {RPULLDOWN}
C_PWM_STUCK_INT PWM_STUCK_INT_NODE GND 1uF
G_PWM_STUCK_INT PWM_STUCK_INT_NODE GND VALUE={V(PWM_STUCK_RAW_NODE)/STUCK_DURATION_THRESHOLD_S}
R_PWM_STUCK_INT_PULLDOWN PWM_STUCK_INT_NODE GND {RPULLDOWN}
E_FAULT_PWM_STUCK FAULT_PWM_STUCK_FLAG GND VALUE={LIMIT(V(PWM_STUCK_INT_NODE)*100, 0, 1)}
R_PWM_STUCK_FLAG_PULLDOWN FAULT_PWM_STUCK_FLAG GND {RPULLDOWN}

* Overtemperature Comparator
E_U10_OVERTEMP FAULT_OVERTEMP_FLAG GND VALUE={MIN(MAX(0.0, (V(TEMP_NODE) - V(/TEMP_THRESHHOLD)))*1k, 1)}
R_OVERTEMP_FLAG_PULLDOWN FAULT_OVERTEMP_FLAG GND {RPULLDOWN}

* Insulation Damage Detection
E_INS_STRESS INS_STRESS_RAW_NODE GND VALUE={V(TEMP_NODE) - 60}
R_INS_STRESS_RAW_PULLDOWN INS_STRESS_RAW_NODE GND {RPULLDOWN}
E_INS_STRESS_NODE INS_STRESS_NODE GND VALUE={MAX(0.0, V(INS_STRESS_RAW_NODE))}
R_INS_STRESS_NODE_PULLDOWN INS_STRESS_NODE GND {RPULLDOWN}
C_INS INT_NODE GND 1u
G_INS INT_NODE GND VALUE={V(INS_STRESS_NODE)/100}
R_INS_INT_NODE_PULLDOWN INT_NODE GND {RPULLDOWN}
E_INS_HEALTH INS_HEALTH_NODE GND VALUE={1 - V(INT_NODE)}
R_INS_HEALTH_PULLDOWN INS_HEALTH_NODE GND {RPULLDOWN}
E_INS_COMP_DIFF FAULT_INS_DIFF_NODE GND VALUE={V(INSULATION_THRESHOLD_NODE) - V(INS_HEALTH_NODE)}
R_INS_COMP_DIFF_PULLDOWN FAULT_INS_DIFF_NODE GND {RPULLDOWN}
E_INS_COMP FAULT_INSULATION_DAMAGE_FLAG GND VALUE={LIMIT(V(FAULT_INS_DIFF_NODE) * 1k, 0, 1)}
R_INS_FLAG_PULLDOWN FAULT_INSULATION_DAMAGE_FLAG GND {RPULLDOWN}

* Sensor Failure Detection
E_SPD_STATIC_ABS SPD_STATIC_ABS_NODE GND VALUE={abs(ddt(V(/MOTOR_SPEED_NODE)))}
R_SPD_STATIC_ABS_PULLDOWN SPD_STATIC_ABS_NODE GND {RPULLDOWN}
E_SPD_STATIC_COND SPD_STATIC_COND_NODE GND VALUE={MIN(MAX(0.0, (0.01 - V(SPD_STATIC_ABS_NODE)))*1k, 1)} ; If ddt is less than 0.01
R_SPD_STATIC_COND_PULLDOWN SPD_STATIC_COND_NODE GND {RPULLDOWN}
E_TIME_COND TIME_COND_NODE GND VALUE={MIN(MAX(0.0, (time - 10u))*1k, 1)} ; If time > 10u
R_TIME_COND_PULLDOWN TIME_COND_NODE GND {RPULLDOWN}
E_SPD_STATIC FAULT_SENSOR_FLAG_RAW GND VALUE={V(SPD_STATIC_COND_NODE) * V(TIME_COND_NODE)}
R_FAULT_SENSOR_RAW_PULLDOWN FAULT_SENSOR_FLAG_RAW GND {RPULLDOWN}
C_SENS SENSOR_INT GND 1u
G_SENS SENSOR_INT GND VALUE={V(FAULT_SENSOR_FLAG_RAW)/STUCK_DURATION_THRESHOLD_S}
R_SENS_INT_PULLDOWN SENSOR_INT GND {RPULLDOWN}
E_SENSOR FAULT_SENSOR_FLAG GND VALUE={LIMIT(V(SENSOR_INT)*100, 0, 1)}
R_SENSOR_FLAG_PULLDOWN FAULT_SENSOR_FLAG GND {RPULLDOWN}

* --- Fault Combination Logic (Behavioral) ---
E_MASTER_FAULT_SUM MASTER_FAULT_SUM_NODE GND VALUE={V(FAULT_OVERCURRENT_FLAG) + V(FAULT_PWM_STUCK_FLAG) + V(FAULT_STALL_FLAG) + V(FAULT_OVERTEMP_FLAG) + V(FAULT_INSULATION_DAMAGE_FLAG) + V(FAULT_SENSOR_FLAG)}
R_MASTER_SUM_PULLDOWN MASTER_FAULT_SUM_NODE GND {RPULLDOWN}
E_MASTER_FAULT MASTER_TRACTION_FAULT GND VALUE={LIMIT(V(MASTER_FAULT_SUM_NODE), 0, 1)}
R_MASTER_FAULT_PULLDOWN MASTER_TRACTION_FAULT GND {RPULLDOWN}

* --- TEG Circuit (KiCAD E2, R10) ---
E2_TEG_OUTPUT Net-_E2-N+_ GND TEMP_NODE GND {TEG_GAIN_VAL}
R10_TEG_LOAD Net-_E2-N+_ GND 100
R_TEG_OUT_PULLDOWN Net-_E2-N+_ GND {RPULLDOWN}

* --- Fault Response / Braking & Regenerative Path ---

* Control signal for braking
E_BRAKE_CTRL_SUM BRAKE_CTRL_SUM_NODE GND VALUE={V(/USER_CONTROLLED_BRAKE) + V(MASTER_TRACTION_FAULT)}
R_BRAKE_CTRL_SUM_PULLDOWN BRAKE_CTRL_SUM_NODE GND {RPULLDOWN}
E_BRAKE_CTRL USER_BRAKE_OR_FAULT_CTRL GND VALUE={LIMIT(V(BRAKE_CTRL_SUM_NODE), 0, 1)}
R_USER_BRAKE_CTRL_PULLDOWN USER_BRAKE_OR_FAULT_CTRL GND {RPULLDOWN}

* Braking Resistor Path (M_BRAKE_RESISTOR, R_BRAKE_RESISTOR) - Parallel to Motor Input
M_BRAKE_RESISTOR MOTOR_RA_LA_NODE USER_BRAKE_OR_FAULT_CTRL BRAKE_RES_SWITCHED_NODE BRAKE_RES_SWITCHED_NODE M_BRAKE_VDMOS
R_BRAKE_RESISTOR BRAKE_RES_SWITCHED_NODE GND {BRAKE_RESISTOR_VAL}

* Regenerative Braking Path (Boost Converter Topology for Charging C_REGEN_MAIN)
L_REGEN_BOOST MOTOR_RA_LA_NODE REGEN_BOOST_SWITCH_NODE {L_REGEN_VAL} ; Inductor in series with motor output (from motor side)
R_L_REGEN_BOOST_DAMP REGEN_BOOST_SWITCH_NODE_DAMP REGEN_BOOST_SWITCH_NODE 1u ; Small series R for inductor DC stability
M_REGEN_BOOST_SWITCH REGEN_BOOST_SWITCH_NODE_DAMP REGEN_CTRL_SIGNAL GND GND __Q3 ; Boost switch (KiCAD Q3 equivalent)
R_REGEN_CTRL_PULLDOWN REGEN_CTRL_SIGNAL GND {RPULLDOWN}
D_REGEN_BOOST_DIODE POWER_DISTRIBUTION_NODE REGEN_BOOST_SWITCH_NODE_DAMP __D1 ; Diode to push current to POWER_DISTRIBUTION_NODE
C_REGEN_MAIN POWER_DISTRIBUTION_NODE GND {REGEN_CAP_VAL} ; Main Regenerative Storage Cap (KiCAD C3 equivalent)
R_C_REGEN_MAIN_SHUNT POWER_DISTRIBUTION_NODE GND 1G ; Shunt across capacitor for DC stability

E_REGEN_CTRL_COND_A REGEN_CTRL_COND_A_NODE GND VALUE={LIMIT((V(/MOTOR_SPEED_NODE) - V(/V_REF)) * 1k, 0, 1)}
R_REGEN_A_PULLDOWN REGEN_CTRL_COND_A_NODE GND {RPULLDOWN}
E_REGEN_CTRL_COND_B REGEN_CTRL_COND_B_NODE GND VALUE={(V(/V_REF) > 0.1 ? 1 : 0)}
R_REGEN_B_PULLDOWN REGEN_CTRL_COND_B_NODE GND {RPULLDOWN}
E_REGEN_CTRL_COND_C REGEN_CTRL_COND_C_NODE GND VALUE={(V(MASTER_TRACTION_FAULT) > 0.5 ? 0 : 1)}
R_REGEN_C_PULLDOWN REGEN_CTRL_COND_C_NODE GND {RPULLDOWN}
E_REGEN_CTRL_SIGNAL REGEN_CTRL_SIGNAL GND VALUE={V(REGEN_CTRL_COND_A_NODE) * V(REGEN_CTRL_COND_B_NODE) * V(REGEN_CTRL_COND_C_NODE)}
R_REGEN_SIGNAL_PULLDOWN REGEN_CTRL_SIGNAL GND {RPULLDOWN}

* --- Temperature Source (Behavioral) ---
E_TEMP_SOURCE TEMP_NODE GND VALUE={25 + (V(CURRENT_SENSE_OUT)*V(CURRENT_SENSE_OUT)*10)}
R_TEMP_NODE_PULLDOWN TEMP_NODE GND {RPULLDOWN}

* --- Simulation Control ---
.control
tran 100u 10s
plot V(/MOTOR_SPEED_NODE) V(/V_REF)
plot V(CURRENT_SENSE_OUT)
plot V(TEMP_NODE)
plot V(MASTER_TRACTION_FAULT)
plot V(PWM_OUT_NODE) V(PID_OUT_NODE)
.endc

.end